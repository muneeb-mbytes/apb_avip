//-------------------------------------------------------
//
//Add HVL_TOP
//-------------------------------------------------------
