//--------------------------------------------------------------------------------------------
// Add Base_test
//--------------------------------------------------------------------------------------------
