//-------------------------------------------------------
//
//Add Slave Driver Bfm
//-------------------------------------------------------
