//-------------------------------------------------------
//
//Add ENV
//-------------------------------------------------------
