//--------------------------------------------------------------------------------------------
// Add APB Virtual Seq PKg
//--------------------------------------------------------------------------------------------
