//-------------------------------------------------------
// Add Slave Agent
//-------------------------------------------------------
