//-------------------------------------------------------
//
//Please Add gloabal Pcakages
//-------------------------------------------------------
