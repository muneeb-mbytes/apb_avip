//-------------------------------------------------------
//
//Add Master Driver Bfm
//-------------------------------------------------------
