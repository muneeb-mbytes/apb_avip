//-------------------------------------------------------
//
//Add Slave Agent Bfm
//-------------------------------------------------------
