//-------------------------------------------------------
//
//Add Master Monitor Bfm
//-------------------------------------------------------
