//-------------------------------------------------------
//
//Add Slave Monitor Bfm
//-------------------------------------------------------
