//-------------------------------------------------------
// Add HDL Top
//-------------------------------------------------------
