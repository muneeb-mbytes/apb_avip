//-------------------------------------------------------
// Add Virtual Sequencer
//-------------------------------------------------------
