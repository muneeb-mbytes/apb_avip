//-------------------------------------------------------
// Add Master Agent 
//-------------------------------------------------------
