//-------------------------------------------------------
//
//Add Master Agent Bfm
//-------------------------------------------------------
