//--------------------------------------------------------------------------------------------
// Slave Base seq
//--------------------------------------------------------------------------------------------
