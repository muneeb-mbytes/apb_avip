//--------------------------------------------------------------------------------------------
// Master Base Seq
//--------------------------------------------------------------------------------------------
