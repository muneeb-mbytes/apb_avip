//-------------------------------------------------------
//Add apb interface 
//-------------------------------------------------------
